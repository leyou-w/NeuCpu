// 6-64译码器模块：将6位输入编码转换为64位独热码输出
// 在CPU设计中用于更广泛的寄存器选择、控制信号生成等场景
// 例如：用于64位寄存器堆的寄存器选择或更复杂的控制信号解码
`include "defines.vh"
module decoder_6_64 (
    input wire [5:0] in,        // 6位输入编码（0-63）
    output reg [63:0] out      // 64位独热码输出（只有1位为1）
);
    // 组合逻辑：根据输入值生成对应的独热码输出
    // 独热码：只有一位为1，其余位为0的二进制编码
    always @ (*) begin
        case(in)
            6'd00:begin out=64'b0000000000000000000000000000000000000000000000000000000000000001; end  // 输入0，输出第0位为1
            6'd01:begin out=64'b0000000000000000000000000000000000000000000000000000000000000010; end  // 输入1，输出第1位为1
            6'd02:begin out=64'b0000000000000000000000000000000000000000000000000000000000000100; end  // 输入2，输出第2位为1
            6'd03:begin out=64'b0000000000000000000000000000000000000000000000000000000000001000; end  // 输入3，输出第3位为1
            6'd04:begin out=64'b0000000000000000000000000000000000000000000000000000000000010000; end  // 输入4，输出第4位为1
            6'd05:begin out=64'b0000000000000000000000000000000000000000000000000000000000100000; end  // 输入5，输出第5位为1
            6'd06:begin out=64'b0000000000000000000000000000000000000000000000000000000001000000; end  // 输入6，输出第6位为1
            6'd07:begin out=64'b0000000000000000000000000000000000000000000000000000000010000000; end  // 输入7，输出第7位为1
            6'd08:begin out=64'b0000000000000000000000000000000000000000000000000000000100000000; end  // 输入8，输出第8位为1
            6'd09:begin out=64'b0000000000000000000000000000000000000000000000000000001000000000; end  // 输入9，输出第9位为1
            6'd10:begin out=64'b0000000000000000000000000000000000000000000000000000010000000000; end  // 输入10，输出第10位为1
            6'd11:begin out=64'b0000000000000000000000000000000000000000000000000000100000000000; end  // 输入11，输出第11位为1
            6'd12:begin out=64'b0000000000000000000000000000000000000000000000000001000000000000; end  // 输入12，输出第12位为1
            6'd13:begin out=64'b0000000000000000000000000000000000000000000000000010000000000000; end  // 输入13，输出第13位为1
            6'd14:begin out=64'b0000000000000000000000000000000000000000000000000100000000000000; end  // 输入14，输出第14位为1
            6'd15:begin out=64'b0000000000000000000000000000000000000000000000001000000000000000; end  // 输入15，输出第15位为1
            6'd16:begin out=64'b0000000000000000000000000000000000000000000000010000000000000000; end  // 输入16，输出第16位为1
            6'd17:begin out=64'b0000000000000000000000000000000000000000000000100000000000000000; end  // 输入17，输出第17位为1
            6'd18:begin out=64'b0000000000000000000000000000000000000000000001000000000000000000; end  // 输入18，输出第18位为1
            6'd19:begin out=64'b0000000000000000000000000000000000000000000010000000000000000000; end  // 输入19，输出第19位为1
            6'd20:begin out=64'b0000000000000000000000000000000000000000000100000000000000000000; end  // 输入20，输出第20位为1
            6'd21:begin out=64'b0000000000000000000000000000000000000000001000000000000000000000; end  // 输入21，输出第21位为1
            6'd22:begin out=64'b0000000000000000000000000000000000000000010000000000000000000000; end  // 输入22，输出第22位为1
            6'd23:begin out=64'b0000000000000000000000000000000000000000100000000000000000000000; end  // 输入23，输出第23位为1
            6'd24:begin out=64'b0000000000000000000000000000000000000001000000000000000000000000; end  // 输入24，输出第24位为1
            6'd25:begin out=64'b0000000000000000000000000000000000000010000000000000000000000000; end  // 输入25，输出第25位为1
            6'd26:begin out=64'b0000000000000000000000000000000000000100000000000000000000000000; end  // 输入26，输出第26位为1
            6'd27:begin out=64'b0000000000000000000000000000000000001000000000000000000000000000; end  // 输入27，输出第27位为1
            6'd28:begin out=64'b0000000000000000000000000000000000010000000000000000000000000000; end  // 输入28，输出第28位为1
            6'd29:begin out=64'b0000000000000000000000000000000000100000000000000000000000000000; end  // 输入29，输出第29位为1
            6'd30:begin out=64'b0000000000000000000000000000000001000000000000000000000000000000; end  // 输入30，输出第30位为1
            6'd31:begin out=64'b0000000000000000000000000000000010000000000000000000000000000000; end  // 输入31，输出第31位为1
            6'd32:begin out=64'b0000000000000000000000000000000100000000000000000000000000000000; end  // 输入32，输出第32位为1
            6'd33:begin out=64'b0000000000000000000000000000001000000000000000000000000000000000; end  // 输入33，输出第33位为1
            6'd34:begin out=64'b0000000000000000000000000000010000000000000000000000000000000000; end  // 输入34，输出第34位为1
            6'd35:begin out=64'b0000000000000000000000000000100000000000000000000000000000000000; end  // 输入35，输出第35位为1
            6'd36:begin out=64'b0000000000000000000000000001000000000000000000000000000000000000; end  // 输入36，输出第36位为1
            6'd37:begin out=64'b0000000000000000000000000010000000000000000000000000000000000000; end  // 输入37，输出第37位为1
            6'd38:begin out=64'b0000000000000000000000000100000000000000000000000000000000000000; end  // 输入38，输出第38位为1
            6'd39:begin out=64'b0000000000000000000000001000000000000000000000000000000000000000; end  // 输入39，输出第39位为1
            6'd40:begin out=64'b0000000000000000000000010000000000000000000000000000000000000000; end  // 输入40，输出第40位为1
            6'd41:begin out=64'b0000000000000000000000100000000000000000000000000000000000000000; end  // 输入41，输出第41位为1
            6'd42:begin out=64'b0000000000000000000001000000000000000000000000000000000000000000; end  // 输入42，输出第42位为1
            6'd43:begin out=64'b0000000000000000000010000000000000000000000000000000000000000000; end  // 输入43，输出第43位为1
            6'd44:begin out=64'b0000000000000000000100000000000000000000000000000000000000000000; end  // 输入44，输出第44位为1
            6'd45:begin out=64'b0000000000000000001000000000000000000000000000000000000000000000; end  // 输入45，输出第45位为1
            6'd46:begin out=64'b0000000000000000010000000000000000000000000000000000000000000000; end  // 输入46，输出第46位为1
            6'd47:begin out=64'b0000000000000000100000000000000000000000000000000000000000000000; end  // 输入47，输出第47位为1
            6'd48:begin out=64'b0000000000000001000000000000000000000000000000000000000000000000; end  // 输入48，输出第48位为1
            6'd49:begin out=64'b0000000000000010000000000000000000000000000000000000000000000000; end  // 输入49，输出第49位为1
            6'd50:begin out=64'b0000000000000100000000000000000000000000000000000000000000000000; end  // 输入50，输出第50位为1
            6'd51:begin out=64'b0000000000001000000000000000000000000000000000000000000000000000; end  // 输入51，输出第51位为1
            6'd52:begin out=64'b0000000000010000000000000000000000000000000000000000000000000000; end  // 输入52，输出第52位为1
            6'd53:begin out=64'b0000000000100000000000000000000000000000000000000000000000000000; end  // 输入53，输出第53位为1
            6'd54:begin out=64'b0000000001000000000000000000000000000000000000000000000000000000; end  // 输入54，输出第54位为1
            6'd55:begin out=64'b0000000010000000000000000000000000000000000000000000000000000000; end  // 输入55，输出第55位为1
            6'd56:begin out=64'b0000000100000000000000000000000000000000000000000000000000000000; end  // 输入56，输出第56位为1
            6'd57:begin out=64'b0000001000000000000000000000000000000000000000000000000000000000; end  // 输入57，输出第57位为1
            6'd58:begin out=64'b0000010000000000000000000000000000000000000000000000000000000000; end  // 输入58，输出第58位为1
            6'd59:begin out=64'b0000100000000000000000000000000000000000000000000000000000000000; end  // 输入59，输出第59位为1
            6'd60:begin out=64'b0001000000000000000000000000000000000000000000000000000000000000; end  // 输入60，输出第60位为1
            6'd61:begin out=64'b0010000000000000000000000000000000000000000000000000000000000000; end  // 输入61，输出第61位为1
            6'd62:begin out=64'b0100000000000000000000000000000000000000000000000000000000000000; end  // 输入62，输出第62位为1
            6'd63:begin out=64'b1000000000000000000000000000000000000000000000000000000000000000; end  // 输入63，输出第63位为1
            default:begin
                out=64'b0;  // 无效输入时输出全0
            end
        endcase
    end

endmodule 