// 5-32译码器模块：将5位输入编码转换为32位独热码输出
// 在CPU设计中用于寄存器选择、控制信号生成等场景
// 例如：将5位寄存器号转换为32位寄存器使能信号
`include "defines.vh"
module decoder_5_32 (
    input wire [4:0] in,        // 5位输入编码（0-31）
    output reg [31:0] out      // 32位独热码输出（只有1位为1）
);
    // 组合逻辑：根据输入值生成对应的独热码输出
    // 独热码：只有一位为1，其余位为0的二进制编码
    always @ (*) begin
        case(in)
            5'd00:begin out=32'b00000000000000000000000000000001; end  // 输入0，输出第0位为1
            5'd01:begin out=32'b00000000000000000000000000000010; end  // 输入1，输出第1位为1
            5'd02:begin out=32'b00000000000000000000000000000100; end  // 输入2，输出第2位为1
            5'd03:begin out=32'b00000000000000000000000000001000; end  // 输入3，输出第3位为1
            5'd04:begin out=32'b00000000000000000000000000010000; end  // 输入4，输出第4位为1
            5'd05:begin out=32'b00000000000000000000000000100000; end  // 输入5，输出第5位为1
            5'd06:begin out=32'b00000000000000000000000001000000; end  // 输入6，输出第6位为1
            5'd07:begin out=32'b00000000000000000000000010000000; end  // 输入7，输出第7位为1
            5'd08:begin out=32'b00000000000000000000000100000000; end  // 输入8，输出第8位为1
            5'd09:begin out=32'b00000000000000000000001000000000; end  // 输入9，输出第9位为1
            5'd10:begin out=32'b00000000000000000000010000000000; end  // 输入10，输出第10位为1
            5'd11:begin out=32'b00000000000000000000100000000000; end  // 输入11，输出第11位为1
            5'd12:begin out=32'b00000000000000000001000000000000; end  // 输入12，输出第12位为1
            5'd13:begin out=32'b00000000000000000010000000000000; end  // 输入13，输出第13位为1
            5'd14:begin out=32'b00000000000000000100000000000000; end  // 输入14，输出第14位为1
            5'd15:begin out=32'b00000000000000001000000000000000; end  // 输入15，输出第15位为1
            5'd16:begin out=32'b00000000000000010000000000000000; end  // 输入16，输出第16位为1
            5'd17:begin out=32'b00000000000000100000000000000000; end  // 输入17，输出第17位为1
            5'd18:begin out=32'b00000000000001000000000000000000; end  // 输入18，输出第18位为1
            5'd19:begin out=32'b00000000000010000000000000000000; end  // 输入19，输出第19位为1
            5'd20:begin out=32'b00000000000100000000000000000000; end  // 输入20，输出第20位为1
            5'd21:begin out=32'b00000000001000000000000000000000; end  // 输入21，输出第21位为1
            5'd22:begin out=32'b00000000010000000000000000000000; end  // 输入22，输出第22位为1
            5'd23:begin out=32'b00000000100000000000000000000000; end  // 输入23，输出第23位为1
            5'd24:begin out=32'b00000001000000000000000000000000; end  // 输入24，输出第24位为1
            5'd25:begin out=32'b00000010000000000000000000000000; end  // 输入25，输出第25位为1
            5'd26:begin out=32'b00000100000000000000000000000000; end  // 输入26，输出第26位为1
            5'd27:begin out=32'b00001000000000000000000000000000; end  // 输入27，输出第27位为1
            5'd28:begin out=32'b00010000000000000000000000000000; end  // 输入28，输出第28位为1
            5'd29:begin out=32'b00100000000000000000000000000000; end  // 输入29，输出第29位为1
            5'd30:begin out=32'b01000000000000000000000000000000; end  // 输入30，输出第30位为1
            5'd31:begin out=32'b10000000000000000000000000000000; end  // 输入31，输出第31位为1
            default:begin
                out=32'b0;  // 无效输入时输出全0
            end
        endcase
    end
endmodule